package Shifter_Ifc;

    import GetPut::*;
    import ClientServer::*;

    typedef Server#(Tuple2#(Bit#(n), Bit #(TLog#(n))), Bit#(n)) Shifter_Ifc #(numeric type n);

endpackage: Shifter_Ifc
